`timescale 1ns / 1ps

////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer:
//
// Create Date:   10:50:05 01/06/2023
// Design Name:   SEQ1011_1007
// Module Name:   C:/Users/admin/Desktop/FPGASDP_120A1107/SEQ1011_1007/SEQ1007_1007_TB.v
// Project Name:  SEQ1011_1007
// Target Device:  
// Tool versions:  
// Description: 
//
// Verilog Test Fixture created by ISE for module: SEQ1011_1007
//
// Dependencies:
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
////////////////////////////////////////////////////////////////////////////////

module SEQ1007_1007_TB;

	// Outputs
	wire ;

	// Instantiate the Unit Under Test (UUT)
	SEQ1011_1007 uut (
		.()
	);

	initial begin
		clk<=0;
		

	end
      
endmodule

